module debug_probe(
    input [31:0] probe_in,
    output [31:0] probe_out
);
    assign probe_out = probe_in;
endmodule 